module pcupdate(
    input clk,
    input [63:0] F_predPC,
    input [63:0] f_valP,f_valC,
    input [3:0]f_icode,
    output reg [63:0] predPC
);

endmodule 